package sine_cordic_constants is

	constant INPUT_DATA_WIDTH    : integer := 8;
    	constant OUTPUT_DATA_WIDTH   : integer := 8;
    	constant ITERATION_COUNT     : integer := 16;
    	constant INTERNAL_PRECISION  : integer := 8;

end sine_cordic_constants;